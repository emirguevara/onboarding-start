module spi_peripheral (
    
);
    
endmodule